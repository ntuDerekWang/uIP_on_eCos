# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Derek Wang
# Original data:  
# Contributors:   
# Date:           2012-4
#
#####DESCRIPTIONEND####
# #uip-udp-packet.c   #uip-ds6.c   tcpip.c    
# ====================================================================
cdl_package CYGPKG_NET_UIP6_STACK {
    display       "uIPv6 Stack"
    description   "ported partially from Contiki uIP Stack"
    hardware
    include_dir   cyg/net/uIPv6Stack/uIPv6
    compile       netstack.c test.c used_sems.c stimer_sys.c timer_sys.c tcpip.c uip6.c uip-udp-packet.c uip-icmp6.c uip-ds6.c random_lib.c list_lib.c ctimer_sys.c uip-debug.c sicslowpan.c packetbuf.c queuebuf.c uip-nd6.c uiplib.c uz2400_dev.c memb_lib.c neighbor-info.c neighbor-attr.c
}
# EOF uIP_stack.cdl
       




