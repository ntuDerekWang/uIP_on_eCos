# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Derek Wang
# Original data:  
# Contributors:   
# Date:           2012-4
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_NET_RIME {
    display       "Rime"
    parent        CYGPKG_NET_UIP6_STACK
    description   "ported partially from Contiki uIP Stack"
    hardware
    include_dir   cyg/net/uIPv6Stack/rime
    compile       rimeaddr.c rimestats.c 
}







